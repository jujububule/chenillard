library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity fonction_2_1 is
port(
    clk_in : in std_logic;
    ledv : buffer std_logic_vector(6 downto 0);
    key2 : in std_logic

);
end fonction_2_1;

architecture chenilleDGDG of fonction_2_1 is

begin
    process(clk_in, key(2))
    begin
        if key2 = '0' then--réinitialisation
				ledv <= "0000000";

			elsif rising_edge(clk_in)then
            case ledv is --permet de décalé la led allumé
                when "0000111" => ledv <= "0001110";
                when "0001110" => ledv <= "0011100";
                when "0011100" => ledv <= "0111000";
                when "0111000" => ledv <= "1110000";
                when "1110000" => ledv <= "0000111";
                when others => ledv <= "0000111";--permet l'initialisation
            end case;
        end if;
    end process;
end chenilleDGDG;
